module teste;
    initial begin
        $display("Icarus Verilog funcionando!");
    end
endmodule